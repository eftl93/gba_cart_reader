module wait_fsm 
						(	input  logic clk,
						input  logic wait_cntr_en,
						input  logic n_reset,
						output logic done
					);
					
					
					
					
					
					
endmodule